module ProcessingBlock(
	input logic [15:0] [15:0] [31:0] initXs,
	input logic [1:0] [15:0] [15:0] [31:0] inWeights,
	input logic [1:0] [15:0] [31:0] inBiases,
	
	
	output logic [16:0] [15:0] [31:0] FinalOut
);

	Processor1 p0(initXs, inWeights, inBiases, FinalOut);
	
	
endmodule