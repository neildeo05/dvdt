/*
 
 VPrime core:
 
 * Contains a 
 
 */



