module Vprime (clk, rst, );

   
endmodule // top
